-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Oct 26 01:06:32 2025


--Name: Phuree Plubjui, Norrapat Kesthong, Vacharavich Ekudomsin
--31 October 2025
--Assignment3

-- Import standard library
LIBRARY ieee;
USE ieee.std_logic_1164.all;

-- Set inputs and outputs
ENTITY FSM_B IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0'; -- active low
        x : IN STD_LOGIC := '0'; --input
        z : OUT STD_LOGIC --output
    );
END FSM_B;

ARCHITECTURE BEHAVIOR OF FSM_B IS
    TYPE type_fstate IS (A,B,C,D,E); -- define finite state machine states
    SIGNAL fstate : type_fstate; -- current state
    SIGNAL reg_fstate : type_fstate; -- next state

BEGIN
---------------------------------------------------------------------
-- Process 1 : State Register
---------------------------------------------------------------------
    PROCESS (clock,reset,reg_fstate)
    BEGIN
        IF (reset='0') THEN -- If reset is active
            fstate <= A; -- go to initial state A
        ELSIF (clock='0' AND clock'event) THEN -- if falling_edge (clock=0)
            fstate <= reg_fstate; -- go to next state
        END IF;
    END PROCESS;

---------------------------------------------------------------------
-- Process 2 : Next State & Output Logic
---------------------------------------------------------------------
    PROCESS (fstate,x)
    BEGIN
        z <= '0';
        CASE fstate IS
		  
				-- State A
            WHEN A =>
                IF (NOT((x = '1'))) THEN -- If x = 0 fo to A
                    reg_fstate <= A;
                ELSIF ((x = '1')) THEN -- If x = 1 fo to B
                    reg_fstate <= B;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= A;
                END IF;

                z <= '0';
					 
				-- State B
            WHEN B =>
                IF (NOT((x = '1'))) THEN -- If x = 0 fo to C
                    reg_fstate <= C;
                ELSIF ((x = '1')) THEN -- If x = 1 fo to B
                    reg_fstate <= B;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= B;
                END IF;

                z <= '0';
					 
				-- State C
            WHEN C =>
                IF (NOT((x = '1'))) THEN -- If x = 0 fo to A
                    reg_fstate <= A;
                ELSIF ((x = '1')) THEN -- If x = 1 fo to D
                    reg_fstate <= D;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= C;
                END IF;

                z <= '0';
					 
				-- State D
            WHEN D =>
                IF (NOT((x = '1'))) THEN -- If x = 0 fo to E
                    reg_fstate <= E;
                ELSIF ((x = '1')) THEN -- If x = 1 fo to B
                    reg_fstate <= B;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= D;
                END IF;

                z <= '0';
				
				-- State E
            WHEN E =>
                IF (NOT((x = '1'))) THEN -- If x = 0 fo to A
                    reg_fstate <= A;
                ELSIF ((x = '1')) THEN -- If x = 1 fo to D
                    reg_fstate <= D;
                -- Inserting 'else' block to prevent latch inference
                ELSE
                    reg_fstate <= E;
                END IF;

                z <= '1';
					 
				-- Default
            WHEN OTHERS => 
                z <= 'X';
                report "Reach undefined state";
        END CASE;
    END PROCESS;
END BEHAVIOR;
